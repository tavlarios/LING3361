BZh91AY&SYˬ� �_�Py���������`	��u+ ��Q�D
BH�
<FBji虑�D�LM���d��6�� MT�j �   2i�# `F&��4� �S!S)6H�D h� � �L�i�����a�0  �@�ѡ�&���F@��M	UR I�|" ��L �5��2		x��$����~wy}/�|+�l�֍!���X�d MK_-e"DA� ��E�.�7�"gt�`τ2��au��b���-⊷K�K�yRKMCI~E���ܷur��z���Ke?����6dx���P4f!�?t��� LA`�$C��-���w�L-fd���T9�<ʵ��y��fk�u���0lRN�{�`�n����[G����%�>�(���I�T���V	3|"�UEJI;cljKAT5�h}�3� U�\@�`1�~����􅘱R!�g<�������'RKJ��t����]fn� ���Zʊd�]]hn;PO�6Օ�h�)r�t3����VӔ{0Dw4@��MMdl<E;u.2�n;B�DcP}�����VoB �lHw:�*X^U%�d����
T!�CTb�2.m����7Y"OC�y�4:��n�w"@.�����=)��� �z�eQV&� ����ԒY)mn2�#R�N�%��Y�9O ��栅Bt�	�xD���pgȼՆ��Y��E�ˈ�	�C&�$�x^H-^���cQ.�bW-b ��)h��KFh<RY;�"v-��z0cm#Q���a�0b�Dz����8ۅ��P��t�HaQ��e���R�Z���K��X�n[�M,V9k��Y��_@g@��1��cm��hi�_��_Yq����zU�2�C6t�����+�I��Ջ%�$��ba"$�j	��)� �B�&40i����J�	�,�	����T�\��0��E�2-j���lBCaV,�Lǔl��p����S���Zo��α0��&��j.���~5�s~��S��f�_墓m�2q��M!!Z���?\Ⱥ�0�y�OC�kő���~���8N��_I�ӻf)� ۜ#��|$���RV_}�G��w%2xD-�\��刀�g�3�$]U���vA�2�[r�z�`���S�:�z���~݃�s�"�*��}$��4A�T�b"J���6)Ϝ����,]e��z�E��iG7*H9��㒾-ӻu��6�l*pɄ�*\|t�"�B�	�1���ހ��w�0zq�B�R�9uT(X�h����"V�AD	�g� Nu�gA�'U�T܌y�kiބ��4�ή����y�ڲUF�ǬB�t��f>���>P������
�@g���-��FY�hs�M�n4�O��������Dd���
h �~]�aUm�KB�&r��CZ{p[�b����M�6D���Bd5�6���`[�Od�}�i������V�0�ؒEݓ� _�^��y�4G�P[ϱ��B��oR�����Q�Q�9��{lU��,�Y$�}�(�V�3M" �6i˔R�T�|�
	�4q���f �bL(T�f�%���f�Ţ�e�k� �H"GA�����s>������	R��C{,�$��ziot{�Tpk�69%3��)D8�b;�r+��8�9¡��@���Fc��E0H��R^aA��$��G���� Ɯ���f�COW4����z��Ea��!0�wsw�j���.�,;�#]�;}�l���;�͕�AE�R(����㽈�$s��������}�01E�ĭ��(UQ�3-w*��3�[�i�r$*BՇ��6"vz5z1Q��B�u>��2�BLa����o@�߁BM�1��۹Q!Z�㼑_�pJ���V���k��:$�3�F��`�ۥb���rE8P�ˬ�